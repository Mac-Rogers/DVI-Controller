`timescale 1ns / 1ps

module main(
    input clk,
    output clk_p,
    output clk_n,
    output red_p,
    output red_n,
    output green_p,
    output green_n,
    output blue_p,
    output blue_n
    );
    
    localparam H_TOTAL = 800;
    localparam V_TOTAL = 525;
    localparam H_ACTIVE = 640;
    localparam V_ACTIVE = 480;
    localparam H_FP = 16; //front porch
    localparam H_BP = 48; //back porch
    localparam V_FP = 10;
    localparam V_BP = 33;
    localparam PINK = 24'hEA63FF;
    localparam GREEN = 24'h5AFF3D;    

    reg pix_clk = 0;
    reg [9:0] hcount = 0;
    reg [9:0] vcount = 0;
    reg [2:0] clk_counter = 0;
    reg hSync, vSync, active_flag;
    reg [23:0] display  = PINK;
    reg [23:0] image_data [1199:0];
    
    // denotes being in the active region
    always @(posedge pix_clk) active_flag <= (hcount < H_ACTIVE) && (vcount < V_ACTIVE);

    // assign sync signals
    always @(posedge pix_clk) hSync <= (hcount > H_ACTIVE + H_FP) && (hcount < H_TOTAL - H_BP);
    always @(posedge pix_clk) vSync <= (vcount > V_ACTIVE + V_FP) && (vcount < V_TOTAL - V_BP);
    
    // assign colours to pattern
    //always @(posedge pix_clk) display <= hcount[6] ? PINK : GREEN;
    always @(posedge pix_clk) display <= image_data[hcount[9:4] + 40*vcount[9:4]];
    
    // creates 10:1 clk divider for 25Mhz
    always @(posedge clk) begin
        if (clk_counter == 4) begin
            clk_counter <= 1'b0;
            pix_clk <= ~pix_clk;
        end else clk_counter <= clk_counter + 1;
    end
    
    // scrolls through grid
    always @(posedge pix_clk) begin
        if (hcount == H_TOTAL) begin
            hcount <= 0; //reset hcount
            vcount <= (vcount == V_TOTAL) ? 1'b0 : vcount + 1; //reset or increment vcount
        end else hcount <= hcount + 1;
    end
    
    // instanciate the encoders
    wire [9:0] TMDS_red, TMDS_green, TMDS_blue;
    TMDS_encoder red_encode(pix_clk, display[23:16], 2'b00, active_flag, TMDS_red);
    TMDS_encoder green_encode(pix_clk, display[15:8], 2'b00, active_flag, TMDS_green);
    TMDS_encoder blue_encode(pix_clk, display[7:0], {vSync,hSync}, active_flag, TMDS_blue);
    
    //serialise the register values
    reg [3:0] TMDS_mod10=0;  // modulus 10 counter
    reg [9:0] TMDS_shift_red=0, TMDS_shift_green=0, TMDS_shift_blue=0;
    reg TMDS_shift_load=0;
    always @(posedge clk) TMDS_shift_load <= (TMDS_mod10==4'd9);

    always @(posedge clk)
    begin
        TMDS_shift_red   <= TMDS_shift_load ? TMDS_red   : TMDS_shift_red  [9:1];
        TMDS_shift_green <= TMDS_shift_load ? TMDS_green : TMDS_shift_green[9:1];
        TMDS_shift_blue  <= TMDS_shift_load ? TMDS_blue  : TMDS_shift_blue [9:1];	
        TMDS_mod10 <= (TMDS_mod10==4'd9) ? 4'd0 : TMDS_mod10+4'd1;
    end
    
    // use the output buffer DS primative to convert single ended signals to diff
    OBUFDS OBUFDS_red  (.I(TMDS_shift_red),   .O(red_p),   .OB(red_n));
    OBUFDS OBUFDS_green(.I(TMDS_shift_green), .O(green_p), .OB(green_n));
    OBUFDS OBUFDS_blue (.I(TMDS_shift_blue),  .O(blue_p),  .OB(blue_n));
    OBUFDS OBUFDS_clk (.I(pix_clk), .O(clk_p), .OB(clk_n));

    initial begin
        image_data[0] = 24'h000000;
        image_data[1] = 24'h000000;
        image_data[2] = 24'h000000;
        image_data[3] = 24'h000000;
        image_data[4] = 24'h000000;
        image_data[5] = 24'h000000;
        image_data[6] = 24'h000000;
        image_data[7] = 24'h000000;
        image_data[8] = 24'h000000;
        image_data[9] = 24'h000000;
        image_data[10] = 24'h000000;
        image_data[11] = 24'h000000;
        image_data[12] = 24'h000000;
        image_data[13] = 24'h000000;
        image_data[14] = 24'h000000;
        image_data[15] = 24'h000000;
        image_data[16] = 24'h000000;
        image_data[17] = 24'h000000;
        image_data[18] = 24'h000000;
        image_data[19] = 24'h000000;
        image_data[20] = 24'h000000;
        image_data[21] = 24'h000000;
        image_data[22] = 24'h000000;
        image_data[23] = 24'h000000;
        image_data[24] = 24'h000000;
        image_data[25] = 24'h000000;
        image_data[26] = 24'h000000;
        image_data[27] = 24'h000000;
        image_data[28] = 24'h000000;
        image_data[29] = 24'h000000;
        image_data[30] = 24'h000000;
        image_data[31] = 24'h000000;
        image_data[32] = 24'h000000;
        image_data[33] = 24'h000000;
        image_data[34] = 24'h000000;
        image_data[35] = 24'h000000;
        image_data[36] = 24'h000000;
        image_data[37] = 24'h000000;
        image_data[38] = 24'h000000;
        image_data[39] = 24'h000000;
        image_data[40] = 24'h000000;
        image_data[41] = 24'h000000;
        image_data[42] = 24'h000000;
        image_data[43] = 24'h000000;
        image_data[44] = 24'h000000;
        image_data[45] = 24'h000000;
        image_data[46] = 24'h000000;
        image_data[47] = 24'h000000;
        image_data[48] = 24'h000000;
        image_data[49] = 24'h000000;
        image_data[50] = 24'h000000;
        image_data[51] = 24'h000000;
        image_data[52] = 24'h000000;
        image_data[53] = 24'h000000;
        image_data[54] = 24'h000000;
        image_data[55] = 24'h000000;
        image_data[56] = 24'h000000;
        image_data[57] = 24'h000000;
        image_data[58] = 24'h000000;
        image_data[59] = 24'h000000;
        image_data[60] = 24'h000000;
        image_data[61] = 24'h000000;
        image_data[62] = 24'h000000;
        image_data[63] = 24'h000000;
        image_data[64] = 24'h000000;
        image_data[65] = 24'h000000;
        image_data[66] = 24'h000000;
        image_data[67] = 24'h000000;
        image_data[68] = 24'h000000;
        image_data[69] = 24'h000000;
        image_data[70] = 24'h000000;
        image_data[71] = 24'h000000;
        image_data[72] = 24'h000000;
        image_data[73] = 24'h000000;
        image_data[74] = 24'h000000;
        image_data[75] = 24'h000000;
        image_data[76] = 24'h000000;
        image_data[77] = 24'h000000;
        image_data[78] = 24'h000000;
        image_data[79] = 24'h000000;
        image_data[80] = 24'h000000;
        image_data[81] = 24'h000000;
        image_data[82] = 24'h000000;
        image_data[83] = 24'h000000;
        image_data[84] = 24'h000000;
        image_data[85] = 24'h000000;
        image_data[86] = 24'h000000;
        image_data[87] = 24'h000000;
        image_data[88] = 24'h000000;
        image_data[89] = 24'h000000;
        image_data[90] = 24'h000000;
        image_data[91] = 24'h000000;
        image_data[92] = 24'h000000;
        image_data[93] = 24'h000000;
        image_data[94] = 24'h000000;
        image_data[95] = 24'h000000;
        image_data[96] = 24'h000000;
        image_data[97] = 24'h000000;
        image_data[98] = 24'h000000;
        image_data[99] = 24'h000000;
        image_data[100] = 24'h000000;
        image_data[101] = 24'h000000;
        image_data[102] = 24'h000000;
        image_data[103] = 24'h000000;
        image_data[104] = 24'h000000;
        image_data[105] = 24'h000000;
        image_data[106] = 24'h000000;
        image_data[107] = 24'h000000;
        image_data[108] = 24'h000000;
        image_data[109] = 24'h000000;
        image_data[110] = 24'h000000;
        image_data[111] = 24'h000000;
        image_data[112] = 24'h000000;
        image_data[113] = 24'h000000;
        image_data[114] = 24'h000000;
        image_data[115] = 24'h000000;
        image_data[116] = 24'h000000;
        image_data[117] = 24'h000000;
        image_data[118] = 24'h000000;
        image_data[119] = 24'h000000;
        image_data[120] = 24'h000000;
        image_data[121] = 24'h000000;
        image_data[122] = 24'h000000;
        image_data[123] = 24'h000000;
        image_data[124] = 24'h000000;
        image_data[125] = 24'h000000;
        image_data[126] = 24'h000000;
        image_data[127] = 24'h000000;
        image_data[128] = 24'h000000;
        image_data[129] = 24'h000000;
        image_data[130] = 24'h000000;
        image_data[131] = 24'h000000;
        image_data[132] = 24'h000000;
        image_data[133] = 24'h000000;
        image_data[134] = 24'h000000;
        image_data[135] = 24'h000000;
        image_data[136] = 24'h000000;
        image_data[137] = 24'h000000;
        image_data[138] = 24'h000000;
        image_data[139] = 24'h000000;
        image_data[140] = 24'h000000;
        image_data[141] = 24'h000000;
        image_data[142] = 24'h000000;
        image_data[143] = 24'h000000;
        image_data[144] = 24'h000000;
        image_data[145] = 24'h000000;
        image_data[146] = 24'h000000;
        image_data[147] = 24'h000000;
        image_data[148] = 24'h000000;
        image_data[149] = 24'h000000;
        image_data[150] = 24'h000000;
        image_data[151] = 24'h000000;
        image_data[152] = 24'h000000;
        image_data[153] = 24'h000000;
        image_data[154] = 24'h000000;
        image_data[155] = 24'h000000;
        image_data[156] = 24'h000000;
        image_data[157] = 24'h000000;
        image_data[158] = 24'h000000;
        image_data[159] = 24'h000000;
        image_data[160] = 24'h000000;
        image_data[161] = 24'h000000;
        image_data[162] = 24'h000000;
        image_data[163] = 24'h000000;
        image_data[164] = 24'h000000;
        image_data[165] = 24'h000000;
        image_data[166] = 24'h000000;
        image_data[167] = 24'h000000;
        image_data[168] = 24'h000000;
        image_data[169] = 24'h000000;
        image_data[170] = 24'h000000;
        image_data[171] = 24'h000000;
        image_data[172] = 24'h000000;
        image_data[173] = 24'h000000;
        image_data[174] = 24'h000000;
        image_data[175] = 24'h000000;
        image_data[176] = 24'h000000;
        image_data[177] = 24'h000000;
        image_data[178] = 24'h000000;
        image_data[179] = 24'h000000;
        image_data[180] = 24'h000000;
        image_data[181] = 24'h000000;
        image_data[182] = 24'h000000;
        image_data[183] = 24'h000000;
        image_data[184] = 24'h000000;
        image_data[185] = 24'h000000;
        image_data[186] = 24'h000000;
        image_data[187] = 24'h000000;
        image_data[188] = 24'h000000;
        image_data[189] = 24'h000000;
        image_data[190] = 24'h000000;
        image_data[191] = 24'h000000;
        image_data[192] = 24'h000000;
        image_data[193] = 24'h000000;
        image_data[194] = 24'h000000;
        image_data[195] = 24'h000000;
        image_data[196] = 24'h000000;
        image_data[197] = 24'h000000;
        image_data[198] = 24'h000000;
        image_data[199] = 24'h000000;
        image_data[200] = 24'h000000;
        image_data[201] = 24'h000000;
        image_data[202] = 24'h000000;
        image_data[203] = 24'h000000;
        image_data[204] = 24'h000000;
        image_data[205] = 24'h000000;
        image_data[206] = 24'h000000;
        image_data[207] = 24'h000000;
        image_data[208] = 24'h000000;
        image_data[209] = 24'h000000;
        image_data[210] = 24'h000000;
        image_data[211] = 24'h000000;
        image_data[212] = 24'h000000;
        image_data[213] = 24'h000000;
        image_data[214] = 24'h000000;
        image_data[215] = 24'h000000;
        image_data[216] = 24'h000000;
        image_data[217] = 24'h000000;
        image_data[218] = 24'h000000;
        image_data[219] = 24'h000000;
        image_data[220] = 24'h000000;
        image_data[221] = 24'h000000;
        image_data[222] = 24'h000000;
        image_data[223] = 24'h000000;
        image_data[224] = 24'h000000;
        image_data[225] = 24'h000000;
        image_data[226] = 24'h000000;
        image_data[227] = 24'h000000;
        image_data[228] = 24'h000000;
        image_data[229] = 24'h000000;
        image_data[230] = 24'h000000;
        image_data[231] = 24'h000000;
        image_data[232] = 24'h000000;
        image_data[233] = 24'h000000;
        image_data[234] = 24'h000000;
        image_data[235] = 24'h000000;
        image_data[236] = 24'h000000;
        image_data[237] = 24'h000000;
        image_data[238] = 24'h000000;
        image_data[239] = 24'h000000;
        image_data[240] = 24'h000000;
        image_data[241] = 24'h000000;
        image_data[242] = 24'h000000;
        image_data[243] = 24'h000000;
        image_data[244] = 24'h000000;
        image_data[245] = 24'h000000;
        image_data[246] = 24'h000000;
        image_data[247] = 24'h000000;
        image_data[248] = 24'h000000;
        image_data[249] = 24'h000000;
        image_data[250] = 24'h000000;
        image_data[251] = 24'h000000;
        image_data[252] = 24'h000000;
        image_data[253] = 24'h000000;
        image_data[254] = 24'h000000;
        image_data[255] = 24'h000000;
        image_data[256] = 24'h000000;
        image_data[257] = 24'h000000;
        image_data[258] = 24'h000000;
        image_data[259] = 24'h000000;
        image_data[260] = 24'h000000;
        image_data[261] = 24'h000000;
        image_data[262] = 24'h000000;
        image_data[263] = 24'h000000;
        image_data[264] = 24'h000000;
        image_data[265] = 24'h000000;
        image_data[266] = 24'h000000;
        image_data[267] = 24'h000000;
        image_data[268] = 24'h000000;
        image_data[269] = 24'h000000;
        image_data[270] = 24'h000000;
        image_data[271] = 24'h000000;
        image_data[272] = 24'h000000;
        image_data[273] = 24'h000000;
        image_data[274] = 24'h000000;
        image_data[275] = 24'h000000;
        image_data[276] = 24'h000000;
        image_data[277] = 24'h000000;
        image_data[278] = 24'h000000;
        image_data[279] = 24'h000000;
        image_data[280] = 24'h000000;
        image_data[281] = 24'h000000;
        image_data[282] = 24'h000000;
        image_data[283] = 24'h000000;
        image_data[284] = 24'h000000;
        image_data[285] = 24'h000000;
        image_data[286] = 24'h000000;
        image_data[287] = 24'h000000;
        image_data[288] = 24'h000000;
        image_data[289] = 24'h000000;
        image_data[290] = 24'h000000;
        image_data[291] = 24'h000000;
        image_data[292] = 24'h000000;
        image_data[293] = 24'h000000;
        image_data[294] = 24'h000000;
        image_data[295] = 24'h000000;
        image_data[296] = 24'h000000;
        image_data[297] = 24'h000000;
        image_data[298] = 24'h000000;
        image_data[299] = 24'h000000;
        image_data[300] = 24'h000000;
        image_data[301] = 24'h000000;
        image_data[302] = 24'h000000;
        image_data[303] = 24'h000000;
        image_data[304] = 24'h000000;
        image_data[305] = 24'h000000;
        image_data[306] = 24'h000000;
        image_data[307] = 24'h000000;
        image_data[308] = 24'h000000;
        image_data[309] = 24'h000000;
        image_data[310] = 24'h000000;
        image_data[311] = 24'h000000;
        image_data[312] = 24'h000000;
        image_data[313] = 24'h000000;
        image_data[314] = 24'h000000;
        image_data[315] = 24'h000000;
        image_data[316] = 24'h000000;
        image_data[317] = 24'h000000;
        image_data[318] = 24'h000000;
        image_data[319] = 24'h000000;
        image_data[320] = 24'h000000;
        image_data[321] = 24'h000000;
        image_data[322] = 24'h000000;
        image_data[323] = 24'h000000;
        image_data[324] = 24'h000000;
        image_data[325] = 24'h000000;
        image_data[326] = 24'h000000;
        image_data[327] = 24'h000000;
        image_data[328] = 24'h000000;
        image_data[329] = 24'h000000;
        image_data[330] = 24'h000000;
        image_data[331] = 24'h000000;
        image_data[332] = 24'h000000;
        image_data[333] = 24'h000000;
        image_data[334] = 24'h000000;
        image_data[335] = 24'h000000;
        image_data[336] = 24'h000000;
        image_data[337] = 24'h000000;
        image_data[338] = 24'h000000;
        image_data[339] = 24'h000000;
        image_data[340] = 24'h000000;
        image_data[341] = 24'h000000;
        image_data[342] = 24'h000000;
        image_data[343] = 24'h000000;
        image_data[344] = 24'h000000;
        image_data[345] = 24'h000000;
        image_data[346] = 24'h000000;
        image_data[347] = 24'h000000;
        image_data[348] = 24'h000000;
        image_data[349] = 24'h000000;
        image_data[350] = 24'h000000;
        image_data[351] = 24'h000000;
        image_data[352] = 24'h000000;
        image_data[353] = 24'h000000;
        image_data[354] = 24'h000000;
        image_data[355] = 24'h000000;
        image_data[356] = 24'h000000;
        image_data[357] = 24'h000000;
        image_data[358] = 24'h000000;
        image_data[359] = 24'h000000;
        image_data[360] = 24'h000000;
        image_data[361] = 24'h000000;
        image_data[362] = 24'h000000;
        image_data[363] = 24'h000000;
        image_data[364] = 24'h000000;
        image_data[365] = 24'h000000;
        image_data[366] = 24'h000000;
        image_data[367] = 24'h000000;
        image_data[368] = 24'h000000;
        image_data[369] = 24'h000000;
        image_data[370] = 24'h000000;
        image_data[371] = 24'h000000;
        image_data[372] = 24'hfe0000;
        image_data[373] = 24'hfe0000;
        image_data[374] = 24'hfe0000;
        image_data[375] = 24'hfe0000;
        image_data[376] = 24'hfe0000;
        image_data[377] = 24'hfe0000;
        image_data[378] = 24'h000000;
        image_data[379] = 24'h000000;
        image_data[380] = 24'h000000;
        image_data[381] = 24'h000000;
        image_data[382] = 24'h000000;
        image_data[383] = 24'h000000;
        image_data[384] = 24'hfe0000;
        image_data[385] = 24'hfe0000;
        image_data[386] = 24'hfe0000;
        image_data[387] = 24'hfe0000;
        image_data[388] = 24'hfe0000;
        image_data[389] = 24'hfe0000;
        image_data[390] = 24'h000000;
        image_data[391] = 24'h000000;
        image_data[392] = 24'h000000;
        image_data[393] = 24'h000000;
        image_data[394] = 24'h000000;
        image_data[395] = 24'h000000;
        image_data[396] = 24'h000000;
        image_data[397] = 24'h000000;
        image_data[398] = 24'h000000;
        image_data[399] = 24'h000000;
        image_data[400] = 24'h000000;
        image_data[401] = 24'h000000;
        image_data[402] = 24'h000000;
        image_data[403] = 24'h000000;
        image_data[404] = 24'h000000;
        image_data[405] = 24'h000000;
        image_data[406] = 24'h000000;
        image_data[407] = 24'h000000;
        image_data[408] = 24'h000000;
        image_data[409] = 24'h000000;
        image_data[410] = 24'h000000;
        image_data[411] = 24'hfe0000;
        image_data[412] = 24'hfe0000;
        image_data[413] = 24'hfe0000;
        image_data[414] = 24'hfd0000;
        image_data[415] = 24'hfd0000;
        image_data[416] = 24'hfd0000;
        image_data[417] = 24'hfe0000;
        image_data[418] = 24'hfe0000;
        image_data[419] = 24'h000000;
        image_data[420] = 24'h000000;
        image_data[421] = 24'h000000;
        image_data[422] = 24'h000000;
        image_data[423] = 24'hfe0000;
        image_data[424] = 24'hfe0000;
        image_data[425] = 24'hfd0000;
        image_data[426] = 24'hfd0000;
        image_data[427] = 24'hfd0000;
        image_data[428] = 24'hfd0000;
        image_data[429] = 24'hfe0000;
        image_data[430] = 24'hfe0000;
        image_data[431] = 24'h000000;
        image_data[432] = 24'h000000;
        image_data[433] = 24'h000000;
        image_data[434] = 24'h000000;
        image_data[435] = 24'h000000;
        image_data[436] = 24'h000000;
        image_data[437] = 24'h000000;
        image_data[438] = 24'h000000;
        image_data[439] = 24'h000000;
        image_data[440] = 24'h000000;
        image_data[441] = 24'h000000;
        image_data[442] = 24'h000000;
        image_data[443] = 24'h000000;
        image_data[444] = 24'h000000;
        image_data[445] = 24'h000000;
        image_data[446] = 24'h000000;
        image_data[447] = 24'h000000;
        image_data[448] = 24'h000000;
        image_data[449] = 24'h000000;
        image_data[450] = 24'hfe0000;
        image_data[451] = 24'hfe0000;
        image_data[452] = 24'hffffff;
        image_data[453] = 24'hffffff;
        image_data[454] = 24'hfe0000;
        image_data[455] = 24'hfe0000;
        image_data[456] = 24'hfe0000;
        image_data[457] = 24'hfe0000;
        image_data[458] = 24'hfe0000;
        image_data[459] = 24'hfe0000;
        image_data[460] = 24'h000000;
        image_data[461] = 24'h000000;
        image_data[462] = 24'hfe0000;
        image_data[463] = 24'hfe0000;
        image_data[464] = 24'hff0000;
        image_data[465] = 24'hfe0000;
        image_data[466] = 24'hfe0000;
        image_data[467] = 24'hfe0000;
        image_data[468] = 24'hff0000;
        image_data[469] = 24'hfe0000;
        image_data[470] = 24'hfe0000;
        image_data[471] = 24'hfe0000;
        image_data[472] = 24'h000000;
        image_data[473] = 24'h000000;
        image_data[474] = 24'h000000;
        image_data[475] = 24'h000000;
        image_data[476] = 24'h000000;
        image_data[477] = 24'h000000;
        image_data[478] = 24'h000000;
        image_data[479] = 24'h000000;
        image_data[480] = 24'h000000;
        image_data[481] = 24'h000000;
        image_data[482] = 24'h000000;
        image_data[483] = 24'h000000;
        image_data[484] = 24'h000000;
        image_data[485] = 24'h000000;
        image_data[486] = 24'h000000;
        image_data[487] = 24'h000000;
        image_data[488] = 24'h000000;
        image_data[489] = 24'hfe0000;
        image_data[490] = 24'hfe0000;
        image_data[491] = 24'hffffff;
        image_data[492] = 24'hffffff;
        image_data[493] = 24'hfe0000;
        image_data[494] = 24'hfe0000;
        image_data[495] = 24'hfe0000;
        image_data[496] = 24'hfe0000;
        image_data[497] = 24'hfe0000;
        image_data[498] = 24'hff0000;
        image_data[499] = 24'hfe0000;
        image_data[500] = 24'hfe0000;
        image_data[501] = 24'hfe0000;
        image_data[502] = 24'hfe0000;
        image_data[503] = 24'hff0000;
        image_data[504] = 24'hfe0000;
        image_data[505] = 24'hfe0000;
        image_data[506] = 24'hfe0000;
        image_data[507] = 24'hfe0000;
        image_data[508] = 24'hfe0000;
        image_data[509] = 24'hfe0000;
        image_data[510] = 24'hff0000;
        image_data[511] = 24'hfe0000;
        image_data[512] = 24'h000000;
        image_data[513] = 24'h000000;
        image_data[514] = 24'h000000;
        image_data[515] = 24'h000000;
        image_data[516] = 24'h000000;
        image_data[517] = 24'h000000;
        image_data[518] = 24'h000000;
        image_data[519] = 24'h000000;
        image_data[520] = 24'h000000;
        image_data[521] = 24'h000000;
        image_data[522] = 24'h000000;
        image_data[523] = 24'h000000;
        image_data[524] = 24'h000000;
        image_data[525] = 24'h000000;
        image_data[526] = 24'h000000;
        image_data[527] = 24'h000000;
        image_data[528] = 24'h000000;
        image_data[529] = 24'hfe0000;
        image_data[530] = 24'hfe0000;
        image_data[531] = 24'hffffff;
        image_data[532] = 24'hfe0000;
        image_data[533] = 24'hfe0000;
        image_data[534] = 24'hfe0000;
        image_data[535] = 24'hfe0000;
        image_data[536] = 24'hfe0000;
        image_data[537] = 24'hfe0000;
        image_data[538] = 24'hff0000;
        image_data[539] = 24'hfd0000;
        image_data[540] = 24'hfe0000;
        image_data[541] = 24'hfe0000;
        image_data[542] = 24'hfe0000;
        image_data[543] = 24'hff0000;
        image_data[544] = 24'hfe0000;
        image_data[545] = 24'hfe0000;
        image_data[546] = 24'hfe0000;
        image_data[547] = 24'hfe0000;
        image_data[548] = 24'hfe0000;
        image_data[549] = 24'hfe0000;
        image_data[550] = 24'hff0000;
        image_data[551] = 24'hfe0000;
        image_data[552] = 24'h000000;
        image_data[553] = 24'h000000;
        image_data[554] = 24'h000000;
        image_data[555] = 24'h000000;
        image_data[556] = 24'h000000;
        image_data[557] = 24'h000000;
        image_data[558] = 24'h000000;
        image_data[559] = 24'h000000;
        image_data[560] = 24'h000000;
        image_data[561] = 24'h000000;
        image_data[562] = 24'h000000;
        image_data[563] = 24'h000000;
        image_data[564] = 24'h000000;
        image_data[565] = 24'h000000;
        image_data[566] = 24'h000000;
        image_data[567] = 24'h000000;
        image_data[568] = 24'h000000;
        image_data[569] = 24'hfe0000;
        image_data[570] = 24'hfe0000;
        image_data[571] = 24'hfe0000;
        image_data[572] = 24'hfe0000;
        image_data[573] = 24'hfe0000;
        image_data[574] = 24'h000000;
        image_data[575] = 24'h000000;
        image_data[576] = 24'h000000;
        image_data[577] = 24'hfe0000;
        image_data[578] = 24'h000000;
        image_data[579] = 24'h000000;
        image_data[580] = 24'h000000;
        image_data[581] = 24'hff0000;
        image_data[582] = 24'h000000;
        image_data[583] = 24'h000000;
        image_data[584] = 24'h000000;
        image_data[585] = 24'hfe0000;
        image_data[586] = 24'h000000;
        image_data[587] = 24'h000000;
        image_data[588] = 24'h000000;
        image_data[589] = 24'hfe0000;
        image_data[590] = 24'hff0000;
        image_data[591] = 24'hfe0000;
        image_data[592] = 24'h000000;
        image_data[593] = 24'h000000;
        image_data[594] = 24'h000000;
        image_data[595] = 24'h000000;
        image_data[596] = 24'h000000;
        image_data[597] = 24'h000000;
        image_data[598] = 24'h000000;
        image_data[599] = 24'h000000;
        image_data[600] = 24'h000000;
        image_data[601] = 24'h000000;
        image_data[602] = 24'h000000;
        image_data[603] = 24'h000000;
        image_data[604] = 24'h000000;
        image_data[605] = 24'h000000;
        image_data[606] = 24'h000000;
        image_data[607] = 24'h000000;
        image_data[608] = 24'h000000;
        image_data[609] = 24'hfe0000;
        image_data[610] = 24'hfe0000;
        image_data[611] = 24'hfe0000;
        image_data[612] = 24'hfe0000;
        image_data[613] = 24'hfe0000;
        image_data[614] = 24'h000000;
        image_data[615] = 24'hfe0000;
        image_data[616] = 24'hfe0000;
        image_data[617] = 24'hfe0000;
        image_data[618] = 24'h000000;
        image_data[619] = 24'hfe0000;
        image_data[620] = 24'h000000;
        image_data[621] = 24'hfe0000;
        image_data[622] = 24'h000000;
        image_data[623] = 24'hfe0000;
        image_data[624] = 24'hfe0000;
        image_data[625] = 24'hfe0000;
        image_data[626] = 24'h000000;
        image_data[627] = 24'hfe0000;
        image_data[628] = 24'h000000;
        image_data[629] = 24'hfe0000;
        image_data[630] = 24'hff0000;
        image_data[631] = 24'hfe0000;
        image_data[632] = 24'h000000;
        image_data[633] = 24'h000000;
        image_data[634] = 24'h000000;
        image_data[635] = 24'h000000;
        image_data[636] = 24'h000000;
        image_data[637] = 24'h000000;
        image_data[638] = 24'h000000;
        image_data[639] = 24'h000000;
        image_data[640] = 24'h000000;
        image_data[641] = 24'h000000;
        image_data[642] = 24'h000000;
        image_data[643] = 24'h000000;
        image_data[644] = 24'h000000;
        image_data[645] = 24'h000000;
        image_data[646] = 24'h000000;
        image_data[647] = 24'h000000;
        image_data[648] = 24'h000000;
        image_data[649] = 24'hfe0000;
        image_data[650] = 24'hfe0000;
        image_data[651] = 24'hfe0000;
        image_data[652] = 24'hfe0000;
        image_data[653] = 24'hfe0000;
        image_data[654] = 24'h000000;
        image_data[655] = 24'h000000;
        image_data[656] = 24'hfe0000;
        image_data[657] = 24'hfe0101;
        image_data[658] = 24'h000000;
        image_data[659] = 24'h000000;
        image_data[660] = 24'h000000;
        image_data[661] = 24'hfe0000;
        image_data[662] = 24'h000000;
        image_data[663] = 24'hfe0000;
        image_data[664] = 24'h000000;
        image_data[665] = 24'hfe0000;
        image_data[666] = 24'h000000;
        image_data[667] = 24'h000000;
        image_data[668] = 24'h000000;
        image_data[669] = 24'hfe0000;
        image_data[670] = 24'hff0000;
        image_data[671] = 24'hfe0000;
        image_data[672] = 24'h000000;
        image_data[673] = 24'h000000;
        image_data[674] = 24'h000000;
        image_data[675] = 24'h000000;
        image_data[676] = 24'h000000;
        image_data[677] = 24'h000000;
        image_data[678] = 24'h000000;
        image_data[679] = 24'h000000;
        image_data[680] = 24'h000000;
        image_data[681] = 24'h000000;
        image_data[682] = 24'h000000;
        image_data[683] = 24'h000000;
        image_data[684] = 24'h000000;
        image_data[685] = 24'h000000;
        image_data[686] = 24'h000000;
        image_data[687] = 24'h000000;
        image_data[688] = 24'h000000;
        image_data[689] = 24'hfe0000;
        image_data[690] = 24'hfe0000;
        image_data[691] = 24'hfc0000;
        image_data[692] = 24'hfe0000;
        image_data[693] = 24'hfe0000;
        image_data[694] = 24'h000000;
        image_data[695] = 24'hfe0303;
        image_data[696] = 24'hfe0000;
        image_data[697] = 24'hfe0000;
        image_data[698] = 24'h000000;
        image_data[699] = 24'hfe0000;
        image_data[700] = 24'hfe0000;
        image_data[701] = 24'hfe0000;
        image_data[702] = 24'h000000;
        image_data[703] = 24'h000000;
        image_data[704] = 24'h000000;
        image_data[705] = 24'hfe0000;
        image_data[706] = 24'h000000;
        image_data[707] = 24'hfe0000;
        image_data[708] = 24'h000000;
        image_data[709] = 24'hfe0000;
        image_data[710] = 24'hfe0000;
        image_data[711] = 24'hfe0000;
        image_data[712] = 24'h000000;
        image_data[713] = 24'h000000;
        image_data[714] = 24'h000000;
        image_data[715] = 24'h000000;
        image_data[716] = 24'h000000;
        image_data[717] = 24'h000000;
        image_data[718] = 24'h000000;
        image_data[719] = 24'h000000;
        image_data[720] = 24'h000000;
        image_data[721] = 24'h000000;
        image_data[722] = 24'h000000;
        image_data[723] = 24'h000000;
        image_data[724] = 24'h000000;
        image_data[725] = 24'h000000;
        image_data[726] = 24'h000000;
        image_data[727] = 24'h000000;
        image_data[728] = 24'h000000;
        image_data[729] = 24'h000000;
        image_data[730] = 24'hfe0000;
        image_data[731] = 24'hfe0000;
        image_data[732] = 24'hff0000;
        image_data[733] = 24'hff0000;
        image_data[734] = 24'hfe0000;
        image_data[735] = 24'hfe0000;
        image_data[736] = 24'hfe0000;
        image_data[737] = 24'hfe0000;
        image_data[738] = 24'hfe0000;
        image_data[739] = 24'hfe0000;
        image_data[740] = 24'hfe0000;
        image_data[741] = 24'hfe0000;
        image_data[742] = 24'hfe0000;
        image_data[743] = 24'hfe0000;
        image_data[744] = 24'hfe0000;
        image_data[745] = 24'hfe0000;
        image_data[746] = 24'hfe0000;
        image_data[747] = 24'hfe0000;
        image_data[748] = 24'hff0000;
        image_data[749] = 24'hfe0000;
        image_data[750] = 24'hfe0000;
        image_data[751] = 24'h000000;
        image_data[752] = 24'h450000;
        image_data[753] = 24'h000000;
        image_data[754] = 24'h000000;
        image_data[755] = 24'h000000;
        image_data[756] = 24'h000000;
        image_data[757] = 24'h000000;
        image_data[758] = 24'h000000;
        image_data[759] = 24'h000000;
        image_data[760] = 24'h000000;
        image_data[761] = 24'h000000;
        image_data[762] = 24'h000000;
        image_data[763] = 24'h000000;
        image_data[764] = 24'h000000;
        image_data[765] = 24'h000000;
        image_data[766] = 24'h000000;
        image_data[767] = 24'h000000;
        image_data[768] = 24'h000000;
        image_data[769] = 24'h000000;
        image_data[770] = 24'h000000;
        image_data[771] = 24'hfe0000;
        image_data[772] = 24'hfe0000;
        image_data[773] = 24'hf50000;
        image_data[774] = 24'hff0000;
        image_data[775] = 24'hfe0000;
        image_data[776] = 24'hfe0000;
        image_data[777] = 24'hfe0000;
        image_data[778] = 24'hfe0000;
        image_data[779] = 24'hfe0000;
        image_data[780] = 24'hfe0000;
        image_data[781] = 24'hfe0000;
        image_data[782] = 24'hfe0000;
        image_data[783] = 24'hfe0000;
        image_data[784] = 24'hfe0000;
        image_data[785] = 24'hfe0000;
        image_data[786] = 24'hfe0000;
        image_data[787] = 24'hff0000;
        image_data[788] = 24'hfe0000;
        image_data[789] = 24'hfe0000;
        image_data[790] = 24'h000000;
        image_data[791] = 24'h000000;
        image_data[792] = 24'h000000;
        image_data[793] = 24'h000000;
        image_data[794] = 24'h000000;
        image_data[795] = 24'h000000;
        image_data[796] = 24'h000000;
        image_data[797] = 24'h000000;
        image_data[798] = 24'h000000;
        image_data[799] = 24'h000000;
        image_data[800] = 24'h000000;
        image_data[801] = 24'h000000;
        image_data[802] = 24'h000000;
        image_data[803] = 24'h000000;
        image_data[804] = 24'h000000;
        image_data[805] = 24'h000000;
        image_data[806] = 24'h000000;
        image_data[807] = 24'h000000;
        image_data[808] = 24'h000000;
        image_data[809] = 24'h000000;
        image_data[810] = 24'h000000;
        image_data[811] = 24'h000000;
        image_data[812] = 24'hfe0000;
        image_data[813] = 24'hfe0000;
        image_data[814] = 24'hff0000;
        image_data[815] = 24'hfe0000;
        image_data[816] = 24'hfe0000;
        image_data[817] = 24'hfe0000;
        image_data[818] = 24'hfe0000;
        image_data[819] = 24'hfe0000;
        image_data[820] = 24'hfe0000;
        image_data[821] = 24'hfe0000;
        image_data[822] = 24'hfe0000;
        image_data[823] = 24'hfe0000;
        image_data[824] = 24'hfe0000;
        image_data[825] = 24'hfe0000;
        image_data[826] = 24'hff0000;
        image_data[827] = 24'hfe0000;
        image_data[828] = 24'hfe0000;
        image_data[829] = 24'h000000;
        image_data[830] = 24'h280000;
        image_data[831] = 24'h000000;
        image_data[832] = 24'h000000;
        image_data[833] = 24'h000000;
        image_data[834] = 24'h000000;
        image_data[835] = 24'h000000;
        image_data[836] = 24'h000000;
        image_data[837] = 24'h000000;
        image_data[838] = 24'h000000;
        image_data[839] = 24'h000000;
        image_data[840] = 24'h000000;
        image_data[841] = 24'h000000;
        image_data[842] = 24'h000000;
        image_data[843] = 24'h000000;
        image_data[844] = 24'h000000;
        image_data[845] = 24'h000000;
        image_data[846] = 24'h000000;
        image_data[847] = 24'h000000;
        image_data[848] = 24'h000000;
        image_data[849] = 24'h000000;
        image_data[850] = 24'h000000;
        image_data[851] = 24'h000000;
        image_data[852] = 24'h000000;
        image_data[853] = 24'hfe0000;
        image_data[854] = 24'hfe0000;
        image_data[855] = 24'hfb0000;
        image_data[856] = 24'hff0000;
        image_data[857] = 24'hfe0000;
        image_data[858] = 24'hfe0000;
        image_data[859] = 24'hfe0000;
        image_data[860] = 24'hfe0000;
        image_data[861] = 24'hfe0000;
        image_data[862] = 24'hfe0000;
        image_data[863] = 24'hfe0000;
        image_data[864] = 24'hfe0000;
        image_data[865] = 24'hff0000;
        image_data[866] = 24'hfe0000;
        image_data[867] = 24'hfe0000;
        image_data[868] = 24'h000000;
        image_data[869] = 24'h000000;
        image_data[870] = 24'h000000;
        image_data[871] = 24'h000000;
        image_data[872] = 24'h000000;
        image_data[873] = 24'h000000;
        image_data[874] = 24'h000000;
        image_data[875] = 24'h000000;
        image_data[876] = 24'h000000;
        image_data[877] = 24'h000000;
        image_data[878] = 24'h000000;
        image_data[879] = 24'h000000;
        image_data[880] = 24'h000000;
        image_data[881] = 24'h000000;
        image_data[882] = 24'h000000;
        image_data[883] = 24'h000000;
        image_data[884] = 24'h000000;
        image_data[885] = 24'h000000;
        image_data[886] = 24'h000000;
        image_data[887] = 24'h000000;
        image_data[888] = 24'h000000;
        image_data[889] = 24'h000000;
        image_data[890] = 24'h000000;
        image_data[891] = 24'h000000;
        image_data[892] = 24'h000000;
        image_data[893] = 24'h000000;
        image_data[894] = 24'hfe0000;
        image_data[895] = 24'hfe0000;
        image_data[896] = 24'hfb0000;
        image_data[897] = 24'hfe0000;
        image_data[898] = 24'hfe0000;
        image_data[899] = 24'hfe0000;
        image_data[900] = 24'hfe0000;
        image_data[901] = 24'hfe0000;
        image_data[902] = 24'hfe0000;
        image_data[903] = 24'hfe0000;
        image_data[904] = 24'hfe0000;
        image_data[905] = 24'hfe0000;
        image_data[906] = 24'hfe0000;
        image_data[907] = 24'h000000;
        image_data[908] = 24'h000000;
        image_data[909] = 24'h000000;
        image_data[910] = 24'h000000;
        image_data[911] = 24'h000000;
        image_data[912] = 24'h000000;
        image_data[913] = 24'h000000;
        image_data[914] = 24'h000000;
        image_data[915] = 24'h000000;
        image_data[916] = 24'h000000;
        image_data[917] = 24'h000000;
        image_data[918] = 24'h000000;
        image_data[919] = 24'h000000;
        image_data[920] = 24'h000000;
        image_data[921] = 24'h000000;
        image_data[922] = 24'h000000;
        image_data[923] = 24'h000000;
        image_data[924] = 24'h000000;
        image_data[925] = 24'h000000;
        image_data[926] = 24'h000000;
        image_data[927] = 24'h000000;
        image_data[928] = 24'h000000;
        image_data[929] = 24'h000000;
        image_data[930] = 24'h000000;
        image_data[931] = 24'h000000;
        image_data[932] = 24'h000000;
        image_data[933] = 24'h000000;
        image_data[934] = 24'h000000;
        image_data[935] = 24'hfe0000;
        image_data[936] = 24'hfe0000;
        image_data[937] = 24'hfe0000;
        image_data[938] = 24'hff0000;
        image_data[939] = 24'hfe0000;
        image_data[940] = 24'hfe0000;
        image_data[941] = 24'hfe0000;
        image_data[942] = 24'hfe0000;
        image_data[943] = 24'hff0000;
        image_data[944] = 24'hfe0000;
        image_data[945] = 24'hfe0000;
        image_data[946] = 24'h000000;
        image_data[947] = 24'h180000;
        image_data[948] = 24'h000000;
        image_data[949] = 24'h000000;
        image_data[950] = 24'h000000;
        image_data[951] = 24'h000000;
        image_data[952] = 24'h000000;
        image_data[953] = 24'h000000;
        image_data[954] = 24'h000000;
        image_data[955] = 24'h000000;
        image_data[956] = 24'h000000;
        image_data[957] = 24'h000000;
        image_data[958] = 24'h000000;
        image_data[959] = 24'h000000;
        image_data[960] = 24'h000000;
        image_data[961] = 24'h000000;
        image_data[962] = 24'h000000;
        image_data[963] = 24'h000000;
        image_data[964] = 24'h000000;
        image_data[965] = 24'h000000;
        image_data[966] = 24'h000000;
        image_data[967] = 24'h000000;
        image_data[968] = 24'h000000;
        image_data[969] = 24'h000000;
        image_data[970] = 24'h000000;
        image_data[971] = 24'h000000;
        image_data[972] = 24'h000000;
        image_data[973] = 24'h000000;
        image_data[974] = 24'h000000;
        image_data[975] = 24'h000000;
        image_data[976] = 24'hfe0000;
        image_data[977] = 24'hfe0000;
        image_data[978] = 24'hf70000;
        image_data[979] = 24'hff0000;
        image_data[980] = 24'hfe0000;
        image_data[981] = 24'hfe0000;
        image_data[982] = 24'hff0000;
        image_data[983] = 24'hfe0000;
        image_data[984] = 24'hfe0000;
        image_data[985] = 24'h000000;
        image_data[986] = 24'h000000;
        image_data[987] = 24'h000000;
        image_data[988] = 24'h000000;
        image_data[989] = 24'h000000;
        image_data[990] = 24'h000000;
        image_data[991] = 24'h000000;
        image_data[992] = 24'h000000;
        image_data[993] = 24'h000000;
        image_data[994] = 24'h000000;
        image_data[995] = 24'h000000;
        image_data[996] = 24'h000000;
        image_data[997] = 24'h000000;
        image_data[998] = 24'h000000;
        image_data[999] = 24'h000000;
        image_data[1000] = 24'h000000;
        image_data[1001] = 24'h000000;
        image_data[1002] = 24'h000000;
        image_data[1003] = 24'h000000;
        image_data[1004] = 24'h000000;
        image_data[1005] = 24'h000000;
        image_data[1006] = 24'h000000;
        image_data[1007] = 24'h000000;
        image_data[1008] = 24'h000000;
        image_data[1009] = 24'h000000;
        image_data[1010] = 24'h000000;
        image_data[1011] = 24'h000000;
        image_data[1012] = 24'h000000;
        image_data[1013] = 24'h000000;
        image_data[1014] = 24'h000000;
        image_data[1015] = 24'h000000;
        image_data[1016] = 24'h000000;
        image_data[1017] = 24'hfe0000;
        image_data[1018] = 24'hfe0000;
        image_data[1019] = 24'hff0000;
        image_data[1020] = 24'hff0000;
        image_data[1021] = 24'hff0000;
        image_data[1022] = 24'hfe0000;
        image_data[1023] = 24'hfe0000;
        image_data[1024] = 24'h000000;
        image_data[1025] = 24'h290000;
        image_data[1026] = 24'h000000;
        image_data[1027] = 24'h000000;
        image_data[1028] = 24'h000000;
        image_data[1029] = 24'h000000;
        image_data[1030] = 24'h000000;
        image_data[1031] = 24'h000000;
        image_data[1032] = 24'h000000;
        image_data[1033] = 24'h000000;
        image_data[1034] = 24'h000000;
        image_data[1035] = 24'h000000;
        image_data[1036] = 24'h000000;
        image_data[1037] = 24'h000000;
        image_data[1038] = 24'h000000;
        image_data[1039] = 24'h000000;
        image_data[1040] = 24'h000000;
        image_data[1041] = 24'h000000;
        image_data[1042] = 24'h000000;
        image_data[1043] = 24'h000000;
        image_data[1044] = 24'h000000;
        image_data[1045] = 24'h000000;
        image_data[1046] = 24'h000000;
        image_data[1047] = 24'h000000;
        image_data[1048] = 24'h000000;
        image_data[1049] = 24'h000000;
        image_data[1050] = 24'h000000;
        image_data[1051] = 24'h000000;
        image_data[1052] = 24'h000000;
        image_data[1053] = 24'h000000;
        image_data[1054] = 24'h000000;
        image_data[1055] = 24'h000000;
        image_data[1056] = 24'h000000;
        image_data[1057] = 24'h000000;
        image_data[1058] = 24'hfe0000;
        image_data[1059] = 24'hfe0000;
        image_data[1060] = 24'hf80000;
        image_data[1061] = 24'hfe0000;
        image_data[1062] = 24'hfe0000;
        image_data[1063] = 24'h000000;
        image_data[1064] = 24'h000000;
        image_data[1065] = 24'h000000;
        image_data[1066] = 24'h000000;
        image_data[1067] = 24'h000000;
        image_data[1068] = 24'h000000;
        image_data[1069] = 24'h000000;
        image_data[1070] = 24'h000000;
        image_data[1071] = 24'h000000;
        image_data[1072] = 24'h000000;
        image_data[1073] = 24'h000000;
        image_data[1074] = 24'h000000;
        image_data[1075] = 24'h000000;
        image_data[1076] = 24'h000000;
        image_data[1077] = 24'h000000;
        image_data[1078] = 24'h000000;
        image_data[1079] = 24'h000000;
        image_data[1080] = 24'h000000;
        image_data[1081] = 24'h000000;
        image_data[1082] = 24'h000000;
        image_data[1083] = 24'h000000;
        image_data[1084] = 24'h000000;
        image_data[1085] = 24'h000000;
        image_data[1086] = 24'h000000;
        image_data[1087] = 24'h000000;
        image_data[1088] = 24'h000000;
        image_data[1089] = 24'h000000;
        image_data[1090] = 24'h000000;
        image_data[1091] = 24'h000000;
        image_data[1092] = 24'h000000;
        image_data[1093] = 24'h000000;
        image_data[1094] = 24'h000000;
        image_data[1095] = 24'h000000;
        image_data[1096] = 24'h000000;
        image_data[1097] = 24'h000000;
        image_data[1098] = 24'h000000;
        image_data[1099] = 24'hfe0000;
        image_data[1100] = 24'hfe0000;
        image_data[1101] = 24'hfe0000;
        image_data[1102] = 24'h000000;
        image_data[1103] = 24'h000000;
        image_data[1104] = 24'h000000;
        image_data[1105] = 24'h000000;
        image_data[1106] = 24'h000000;
        image_data[1107] = 24'h000000;
        image_data[1108] = 24'h000000;
        image_data[1109] = 24'h000000;
        image_data[1110] = 24'h000000;
        image_data[1111] = 24'h000000;
        image_data[1112] = 24'h000000;
        image_data[1113] = 24'h000000;
        image_data[1114] = 24'h000000;
        image_data[1115] = 24'h000000;
        image_data[1116] = 24'h000000;
        image_data[1117] = 24'h000000;
        image_data[1118] = 24'h000000;
        image_data[1119] = 24'h000000;
        image_data[1120] = 24'h000000;
        image_data[1121] = 24'h000000;
        image_data[1122] = 24'h000000;
        image_data[1123] = 24'h000000;
        image_data[1124] = 24'h000000;
        image_data[1125] = 24'h000000;
        image_data[1126] = 24'h000000;
        image_data[1127] = 24'h000000;
        image_data[1128] = 24'h000000;
        image_data[1129] = 24'h000000;
        image_data[1130] = 24'h000000;
        image_data[1131] = 24'h000000;
        image_data[1132] = 24'h000000;
        image_data[1133] = 24'h000000;
        image_data[1134] = 24'h000000;
        image_data[1135] = 24'h000000;
        image_data[1136] = 24'h000000;
        image_data[1137] = 24'h000000;
        image_data[1138] = 24'h000000;
        image_data[1139] = 24'h000000;
        image_data[1140] = 24'h000000;
        image_data[1141] = 24'h000000;
        image_data[1142] = 24'h000000;
        image_data[1143] = 24'h000000;
        image_data[1144] = 24'h000000;
        image_data[1145] = 24'h000000;
        image_data[1146] = 24'h000000;
        image_data[1147] = 24'h000000;
        image_data[1148] = 24'h000000;
        image_data[1149] = 24'h000000;
        image_data[1150] = 24'h000000;
        image_data[1151] = 24'h000000;
        image_data[1152] = 24'h000000;
        image_data[1153] = 24'h000000;
        image_data[1154] = 24'h000000;
        image_data[1155] = 24'h000000;
        image_data[1156] = 24'h000000;
        image_data[1157] = 24'h000000;
        image_data[1158] = 24'h000000;
        image_data[1159] = 24'h000000;
        image_data[1160] = 24'h000000;
        image_data[1161] = 24'h000000;
        image_data[1162] = 24'h000000;
        image_data[1163] = 24'h000000;
        image_data[1164] = 24'h000000;
        image_data[1165] = 24'h000000;
        image_data[1166] = 24'h000000;
        image_data[1167] = 24'h000000;
        image_data[1168] = 24'h000000;
        image_data[1169] = 24'h000000;
        image_data[1170] = 24'h000000;
        image_data[1171] = 24'h000000;
        image_data[1172] = 24'h000000;
        image_data[1173] = 24'h000000;
        image_data[1174] = 24'h000000;
        image_data[1175] = 24'h000000;
        image_data[1176] = 24'h000000;
        image_data[1177] = 24'h000000;
        image_data[1178] = 24'h000000;
        image_data[1179] = 24'h000000;
        image_data[1180] = 24'h000000;
        image_data[1181] = 24'h000000;
        image_data[1182] = 24'h000000;
        image_data[1183] = 24'h000000;
        image_data[1184] = 24'h000000;
        image_data[1185] = 24'h000000;
        image_data[1186] = 24'h000000;
        image_data[1187] = 24'h000000;
        image_data[1188] = 24'h000000;
        image_data[1189] = 24'h000000;
        image_data[1190] = 24'h000000;
        image_data[1191] = 24'h000000;
        image_data[1192] = 24'h000000;
        image_data[1193] = 24'h000000;
        image_data[1194] = 24'h000000;
        image_data[1195] = 24'h000000;
        image_data[1196] = 24'h000000;
        image_data[1197] = 24'h000000;
        image_data[1198] = 24'h000000;
        image_data[1199] = 24'h000000;
    end

endmodule


